----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:31:58 05/20/2022 
-- Design Name: 
-- Module Name:    MUX_4x1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUX_4x1 is
    Port ( inputA : in  STD_LOGIC_VECTOR (31 downto 0);
           inputB : in 	STD_LOGIC_VECTOR (31 downto 0);
           inputC : in  STD_LOGIC_VECTOR (31 downto 0);
			  inputD : in 	STD_LOGIC_VECTOR (31 downto 0);
           Selector : in  STD_LOGIC_VECTOR (1 downto 0);
           MuxOut : out  STD_LOGIC_VECTOR (31 downto 0));
end MUX_4x1;

architecture Behavioral of MUX_4x1 is

begin
	with Selector select
		MuxOut <= InputA when "00",
					  InputB when "01",
					  InputC when "10",
					  InputD when others;
end Behavioral;

