----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    05:22:55 05/18/2022 
-- Design Name: 
-- Module Name:    GenericRegister - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity GenericRegister is
	 generic ( Size : Integer); --Size we want
	 Port ( CLK : in  STD_LOGIC;
           RST : in  STD_LOGIC;
           WE : in  STD_LOGIC;
           Datain : in  STD_LOGIC_VECTOR (Size - 1 downto 0);
           Dataout : out  STD_LOGIC_VECTOR (Size - 1 downto 0));
end GenericRegister;

architecture Behavioral of GenericRegister is

begin
	process (CLK) is 
	begin 		
		if rising_edge(CLK) then
			if RST = '1' then
				Dataout <= (others => '0') after 10ns;
			elsif WE = '1' then
				Dataout <= Datain after 10ns;
			end if;
		end if;
	end process;
	
end Behavioral;

